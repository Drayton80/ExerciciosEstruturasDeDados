library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use STD.TEXTIO.ALL;

entity testbench_divideby3FSM is
	-- no inputs or outputs
end;

architecture sim of testbench_divideby3FSM is
	component divideby3FSM
		port (clk, reset: in STD_LOGIC;
			  y: out STD_LOGIC);
	end component;

signal clk, reset, y, yexpected: STD_LOGIC;
constant MEMSIZE: integer := 11;
type tvarray is array (MEMSIZE downto 0) of STD_LOGIC_VECTOR (1 downto 0);
signal testvectors: tvarray;
shared variable vectornum, errors: integer;

begin
-- instantiate device under test
dut: divideby3FSM port map (clk, reset, y);
-- generate clock
process begin
	clk <= '1'; wait for 10 ns;  
	clk <= '0'; wait for 10 ns;
end process;
-- at start of test, load vectors
-- and pulse reset
process is
file tv: TEXT;
variable i, j: integer;
variable L: line;
variable ch: character;
begin
	-- read file of test vectors
	i := 0;
	FILE_OPEN (tv, "./example.tv", READ_MODE);
	while not endfile(tv) loop
		readline (tv, L);
		for j in 1 downto 0 loop
			read (L, ch);
			
			if (ch = '0') then
				testvectors (i) (j) <= '0';
			else
				testvectors (i) (j) <= '1';
			end if;
			
		end loop;
		i := i + 1;
	end loop;
	vectornum := 0; errors := 0;
	-- reset <= '1'; wait for 27 ns; reset <= '0';
	wait;
end process;
-- apply test vectors on rising edge of clk
process (clk) begin
	if (clk'event and clk='1') then   
		reset <= testvectors (vectornum) (1);
		yexpected <= testvectors (vectornum)(0);
	end if;
end process;
-- check results on falling edge of clk
process (clk) begin
	if (clk'event and clk = '0')then
		assert y = yexpected
			report "Vetor deu erro n. Teste: " &integer'image(vectornum)&
					 ". Esperado yesp ="& STD_LOGIC'image(yexpected)&
					 "Valor Obtido: y ="& STD_LOGIC'image(y);
			
		if (y /= yexpected) then
			errors := errors + 1;
		end if;
		
		vectornum := vectornum + 1;
		-- if (is_x (testvectors(vectornum))) then
		if (vectornum = MEMSIZE) then
			if (errors = 0) then
				report "Just kidding --" &
				integer'image (vectornum) &
				"tests completed successfully."
				severity failure;
			else
				report integer'image (vectornum) &
				"tests completed, errors = " &
				integer'image (errors)
				severity failure;
			end if;
		end if;
	end if;
	
end process;
end;
